module top_module ( input a, input b, output out );
    mod_a ia(a, b, out);
endmodule
